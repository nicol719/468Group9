// ALU Testbench

//================
//ALU Main Module
//================
// Code here


//==================
// 32-bit adder
//=================
//Code here

//==================
// 32-bit subtractor
//=================
//Code here

//==================
// 32-bit multiplier
//=================
//Code here

//==================
// 32-bit bitwise ORing
//=================
//Code here

//==================
// 32-bit bitwise ANDing
//=================
//Code here

//==================
// 32-bit bitwise XORing
//=================
//Code here

//==================
// parameterized 32-bit right shift register that shifts the input by n-bit
//=================
//Code here

//==================
// parameterized 32-bit left shift register that shifts the input by n-bit
//=================
//Code here

//==================
// parameterized 32-bit register that right rotates the input by n-bit
//=================
//Code here

//==================
// A 32-line 16x1 Multiplexer (each input/output is an 32-bit wide)
//=================
//Code here

//==================
// A module that checks the S-bit /CMP instruction and generates the 4-bit flag accordingly
//=================
//Code here

//==================
// 8-bit Counter (Program Counter (PC))
//=================
//Code here


//================
// Other small modules that cover the remaining functions of the 15-instruction set (such as MOV and LDR).
//================