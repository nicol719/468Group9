// Register Bank Here
// Register Bank consists of a 4 to 16 decoder, 16 32-bit registers, and 2 32-bit 16 x 1 mux's

module register_bank;
	//register bank code here
endmodule

module decoder_4to16;
	//decoder code goes here
endmodule

module register_32bit;
	//register code goes here
endmodule

module mux_16x1;
	//mux code goes here
endmodule